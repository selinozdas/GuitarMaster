`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.12.2016 04:10:02
// Design Name: 
// Module Name: songData
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module songData(input logic clk, [12:0] addr,output logic [9:0] data);
reg [9:0] data;
reg [9:0] notes [0:1199];

initial begin
	// initialize the notes
	notes[0] =  10'b0000000000;
	notes[1] =  10'b0000000000;
	notes[2] =  10'b0000000000;
	notes[3] =  10'b0000000000;
	notes[4] =  10'b0000000000;
	notes[5] =  10'b0000000000;
	notes[6] =  10'b0000000000;
	notes[7] =  10'b0000000000;
	notes[8] =  10'b0000000000;
	notes[9] =  10'b0000000000;
	notes[10] = 10'b0000000000;
	notes[11] = 10'b0000000000;
	notes[12] = 10'b0000000000;
	notes[13] = 10'b0000000000;
	notes[14] = 10'b0000000000;
	notes[15] = 10'b0000000000;
	notes[16] = 10'b0010000100; // measure 5, start of song
	notes[17] = 10'b0010000100;
	notes[18] = 10'b0000000000;
	notes[19] = 10'b0010000100;
	notes[20] = 10'b0001000010;
	notes[21] = 10'b0000000000;
	notes[22] = 10'b0001000010;
	notes[23] = 10'b0000000000;
	notes[24] = 10'b0100001000; // 6
	notes[25] = 10'b0100001000;
	notes[26] = 10'b0000000000;
	notes[27] = 10'b0100001000;
	notes[28] = 10'b0100001000;
	notes[29] = 10'b0100001000;
	notes[30] = 10'b0000000000;
	notes[31] = 10'b0100001000;
	notes[32] = 10'b0010000100; // 7
	notes[33] = 10'b0010000100;
	notes[34] = 10'b0000000000;
	notes[35] = 10'b0010000100;
	notes[36] = 10'b0001000010;
	notes[37] = 10'b0000000000;
	notes[38] = 10'b0001000010;
	notes[39] = 10'b0000000000;
	notes[40] = 10'b1000010000; // 8
	notes[41] = 10'b1000010000;
	notes[42] = 10'b0000000000;
	notes[43] = 10'b1000010000;
	notes[44] = 10'b1000010000;
	notes[45] = 10'b1000010000;
	notes[46] = 10'b0000000000;
	notes[47] = 10'b0000000000;
	notes[48] = 10'b0010000100; // 9
	notes[49] = 10'b0010000100;
	notes[50] = 10'b0000000000;
	notes[51] = 10'b0010000100;
	notes[52] = 10'b0001000010;
	notes[53] = 10'b0000000000;
	notes[54] = 10'b0001000010;
	notes[55] = 10'b0000000000;
	notes[56] = 10'b0100001000; // 10
	notes[57] = 10'b0100001000;
	notes[58] = 10'b0000000000;
	notes[59] = 10'b0100001000;
	notes[60] = 10'b0100001000;
	notes[61] = 10'b0100001000;
	notes[62] = 10'b0000000000;
	notes[63] = 10'b0100001000;
	notes[64] = 10'b0010000100; // 11
	notes[65] = 10'b0010000100;
	notes[66] = 10'b0000000000;
	notes[67] = 10'b0010000100;
	notes[68] = 10'b0001000010;
	notes[69] = 10'b0000000000;
	notes[70] = 10'b0001000010;
	notes[71] = 10'b0000000000;
	notes[72] = 10'b0010010000; // 12
	notes[73] = 10'b0010001000;
	notes[74] = 10'b0010000100;
	notes[75] = 10'b0010000000;
	notes[76] = 10'b0100000100;
	notes[77] = 10'b0100000010;
	notes[78] = 10'b0100000010;
	notes[79] = 10'b0100000000;
	notes[80] = 10'b0010001100; // 13
	notes[81] = 10'b0010001100;
	notes[82] = 10'b0000000000;
	notes[83] = 10'b0010000100;
	notes[84] = 10'b0001000010;
	notes[85] = 10'b0000000000;
	notes[86] = 10'b0001000010;
	notes[87] = 10'b0000000000;
	notes[88] = 10'b0100010100; // 14
	notes[89] = 10'b0100010100;
	notes[90] = 10'b0000000000;
	notes[91] = 10'b0100010100;
	notes[92] = 10'b0100010100;
	notes[93] = 10'b0100010100;
	notes[94] = 10'b0000000000;
	notes[95] = 10'b0100010100;
	notes[96] = 10'b0010001100; // 15
	notes[97] = 10'b0010001100;
	notes[98] = 10'b0000000000;
	notes[99] = 10'b0010000100;
	notes[100] = 10'b0001000010;
	notes[101] = 10'b0000000000;
	notes[102] = 10'b0001000010;
	notes[103] = 10'b0000000000;
	notes[104] = 10'b1000011000; // 16
	notes[105] = 10'b1000011000;
	notes[106] = 10'b0000000000;
	notes[107] = 10'b1000011000;
	notes[108] = 10'b1000011000;
	notes[109] = 10'b1000011000;
	notes[110] = 10'b0000000000;
	notes[111] = 10'b0000011000;
	notes[112] = 10'b0010001100; // 17
	notes[113] = 10'b0010001100;
	notes[114] = 10'b0000000000;
	notes[115] = 10'b0010000100;
	notes[116] = 10'b0001000010;
	notes[117] = 10'b0000000000;
	notes[118] = 10'b0001000010;
	notes[119] = 10'b0000000000;
	notes[120] = 10'b0100010100; // 18
	notes[121] = 10'b0100010100;
	notes[122] = 10'b0000000000;
	notes[123] = 10'b0100010100;
	notes[124] = 10'b0100010100;
	notes[125] = 10'b0100010100;
	notes[126] = 10'b0000000000;
	notes[127] = 10'b0100010100;
	notes[128] = 10'b0010001100; // 19
	notes[129] = 10'b0010001100;
	notes[130] = 10'b0000000000;
	notes[131] = 10'b0010000100;
	notes[132] = 10'b0001000010;
	notes[133] = 10'b0000000000;
	notes[134] = 10'b0001000010;
	notes[135] = 10'b0000000000;
	notes[136] = 10'b0010001010; // 20
	notes[137] = 10'b0010001010;
	notes[138] = 10'b0010001010;
	notes[139] = 10'b0010000000;
	notes[140] = 10'b0100001100;
	notes[141] = 10'b0100001100;
	notes[142] = 10'b0100001100;
	notes[143] = 10'b0000000000;
	notes[144] = 10'b0010001000; // 21
	notes[145] = 10'b0010000000;
	notes[146] = 10'b0000001000;
	notes[147] = 10'b0010001000;
	notes[148] = 10'b0001001000;
	notes[149] = 10'b0000000100;
	notes[150] = 10'b0001001000;
	notes[151] = 10'b0000000100;
	notes[152] = 10'b0100001000; // 22
	notes[153] = 10'b0100000000;
	notes[154] = 10'b0000001000;
	notes[155] = 10'b0100001000;
	notes[156] = 10'b0100001000;
	notes[157] = 10'b0100000100;
	notes[158] = 10'b0000001000;
	notes[159] = 10'b0100000100;
	notes[160] = 10'b0010001000; // 23
	notes[161] = 10'b0010000000;
	notes[162] = 10'b0000001000;
	notes[163] = 10'b0010001000;
	notes[164] = 10'b0001001000;
	notes[165] = 10'b0000000100;
	notes[166] = 10'b0001001000;
	notes[167] = 10'b0000000100;
	notes[168] = 10'b1000001000; // 24
	notes[169] = 10'b1000000000;
	notes[170] = 10'b0000001000;
	notes[171] = 10'b1000001000;
	notes[172] = 10'b1000001000;
	notes[173] = 10'b1000010000;
	notes[174] = 10'b0000010000;
	notes[175] = 10'b0000010000;
	notes[176] = 10'b0010001000; // 25
	notes[177] = 10'b0010000000;
	notes[178] = 10'b0000001000;
	notes[179] = 10'b0010001000;
	notes[180] = 10'b0001001000;
	notes[181] = 10'b0000000100;
	notes[182] = 10'b0001001000;
	notes[183] = 10'b0000000100;
	notes[184] = 10'b0100001000; // 26
	notes[185] = 10'b0100000000;
	notes[186] = 10'b0000001000;
	notes[187] = 10'b0100001000;
	notes[188] = 10'b0100001000;
	notes[189] = 10'b0100000100;
	notes[190] = 10'b0000001000;
	notes[191] = 10'b0100000100;
	notes[192] = 10'b0010001000; // 27
	notes[193] = 10'b0010000000;
	notes[194] = 10'b0000001000;
	notes[195] = 10'b0010001000;
	notes[196] = 10'b0001001000;
	notes[197] = 10'b0000000100;
	notes[198] = 10'b0001001000;
	notes[199] = 10'b0000000100;
	notes[200] = 10'b0010000010; // 28
	notes[201] = 10'b0010000000;
	notes[202] = 10'b0010000010;
	notes[203] = 10'b0010000010;
	notes[204] = 10'b0100000010;
	notes[205] = 10'b0100000001;
	notes[206] = 10'b0100000001;
	notes[207] = 10'b0100000000;
	notes[208] = 10'b0001001010; // 29
	notes[209] = 10'b0001001010;
	notes[210] = 10'b0001001010;
	notes[211] = 10'b0001001010;
	notes[212] = 10'b0001001010;
	notes[213] = 10'b0001001010;
	notes[214] = 10'b0001001010;
	notes[215] = 10'b0001000000;
	notes[216] = 10'b0100010100; // 30
	notes[217] = 10'b0100010100;
	notes[218] = 10'b0100010100;
	notes[219] = 10'b0100010100;
	notes[220] = 10'b0100010100;
	notes[221] = 10'b0000000000;
	notes[222] = 10'b0000000000;
	notes[223] = 10'b0000000000;
	notes[224] = 10'b1000001010; // 31
	notes[225] = 10'b0000000000;
	notes[226] = 10'b1000001010;
	notes[227] = 10'b0000000000;
	notes[228] = 10'b1000001010;
	notes[229] = 10'b0100000000;
	notes[230] = 10'b1000001010;
	notes[231] = 10'b0000000000;
	notes[232] = 10'b0010001100; // 32
	notes[233] = 10'b0000000000;
	notes[234] = 10'b0010001100;
	notes[235] = 10'b0000000000;
	notes[236] = 10'b0010001100;
	notes[237] = 10'b0000100000;
	notes[238] = 10'b0010001100;
	notes[239] = 10'b0000000000;
	notes[240] = 10'b1000010010; // 33
	notes[241] = 10'b0000000000;
	notes[242] = 10'b1000010010;
	notes[243] = 10'b0000000000;
	notes[244] = 10'b1000010010;
	notes[245] = 10'b0010000000;
	notes[246] = 10'b1000010010;
	notes[247] = 10'b0000000000;
	notes[248] = 10'b0100000101; // 34
	notes[249] = 10'b0100000000;
	notes[250] = 10'b0100000101;
	notes[251] = 10'b0100000000;
	notes[252] = 10'b0010000110;
	notes[253] = 10'b0010000000;
	notes[254] = 10'b0010000110;
	notes[255] = 10'b0010000000;
	notes[256] = 10'b0001001010; // 35
	notes[257] = 10'b0000000000;
	notes[258] = 10'b0001001010;
	notes[259] = 10'b0000000000;
	notes[260] = 10'b0001001010;
	notes[261] = 10'b0000100000;
	notes[262] = 10'b0001001010;
	notes[263] = 10'b0000000000;
	notes[264] = 10'b0010001100; // 36
	notes[265] = 10'b0000000000;
	notes[266] = 10'b0010001100;
	notes[267] = 10'b0000000000;
	notes[268] = 10'b0010001100;
	notes[269] = 10'b0001000000;
	notes[270] = 10'b0010001100;
	notes[271] = 10'b0000000000;
	notes[272] = 10'b1000010010; // 37
	notes[273] = 10'b0000000000;
	notes[274] = 10'b1000010010;
	notes[275] = 10'b0000000000;
	notes[276] = 10'b1000010010;
	notes[277] = 10'b0010000000;
	notes[278] = 10'b1000010010;
	notes[279] = 10'b0000000000;
	notes[280] = 10'b0100000101; // 38
	notes[281] = 10'b0100000000;
	notes[282] = 10'b0100000101;
	notes[283] = 10'b0100000000;
	notes[284] = 10'b0010000110;
	notes[285] = 10'b0010000000;
	notes[286] = 10'b0010000110;
	notes[287] = 10'b0010000000;
	notes[288] = 10'b0001001010; // 39
	notes[289] = 10'b0000000000;
	notes[290] = 10'b0001001010;
	notes[291] = 10'b0000000000;
	notes[292] = 10'b0001001010;
	notes[293] = 10'b0000000000;
	notes[294] = 10'b0001001010;
	notes[295] = 10'b0000000000;
	notes[296] = 10'b0001001010; // 40
	notes[297] = 10'b0000000000;
	notes[298] = 10'b0001001010;
	notes[299] = 10'b0000000000;
	notes[300] = 10'b0001001010;
	notes[301] = 10'b0010000101;
	notes[302] = 10'b0010000101;
	notes[303] = 10'b0010000000;
	notes[304] = 10'b1000000110; // 41
	notes[305] = 10'b0000000000;
	notes[306] = 10'b1000000110;
	notes[307] = 10'b0000000000;
	notes[308] = 10'b1000000110;
	notes[309] = 10'b0000000000;
	notes[310] = 10'b1000000110;
	notes[311] = 10'b0000000000;
	notes[312] = 10'b1000000110; // 42
	notes[313] = 10'b0000000000;
	notes[314] = 10'b1000000110;
	notes[315] = 10'b0000000000;
	notes[316] = 10'b1000000110;
	notes[317] = 10'b0100000101;
	notes[318] = 10'b0100000101;
	notes[319] = 10'b0010000000;
	notes[320] = 10'b0001001010; // 43
	notes[321] = 10'b0000000000;
	notes[322] = 10'b0001001010;
	notes[323] = 10'b0000000000;
	notes[324] = 10'b0001001010;
	notes[325] = 10'b0000000000;
	notes[326] = 10'b0001001010;
	notes[327] = 10'b0000000000;
	notes[328] = 10'b0001001010; // 44
	notes[329] = 10'b0000000000;
	notes[330] = 10'b0001001010;
	notes[331] = 10'b0000000000;
	notes[332] = 10'b0001001010;
	notes[333] = 10'b0010000101;
	notes[334] = 10'b0010000101;
	notes[335] = 10'b0010000000;
	notes[336] = 10'b1000000110; // 45
	notes[337] = 10'b0000000000;
	notes[338] = 10'b1000000110;
	notes[339] = 10'b0000000000;
	notes[340] = 10'b1000000110;
	notes[341] = 10'b0000000000;
	notes[342] = 10'b1000000110;
	notes[343] = 10'b0000000000;
	notes[344] = 10'b0010000001; // 46
	notes[345] = 10'b0010000001;
	notes[346] = 10'b0010000001;
	notes[347] = 10'b0010000001;
	notes[348] = 10'b0100000010;
	notes[349] = 10'b0000000000;
	notes[350] = 10'b0000000000;
	notes[351] = 10'b0000000000;
	notes[352] = 10'b0010000100; // 47
	notes[353] = 10'b0010000100;
	notes[354] = 10'b0000000000;
	notes[355] = 10'b0010000100;
	notes[356] = 10'b0001000010;
	notes[357] = 10'b0000000000;
	notes[358] = 10'b0001000010;
	notes[359] = 10'b0000000000;
	notes[360] = 10'b0100001000; // 48
	notes[361] = 10'b0100001000;
	notes[362] = 10'b0000000000;
	notes[363] = 10'b0100001000;
	notes[364] = 10'b0100001000;
	notes[365] = 10'b0100001000;
	notes[366] = 10'b0000000000;
	notes[367] = 10'b0100001000;
	notes[368] = 10'b0010000100; // 49
	notes[369] = 10'b0010000100;
	notes[370] = 10'b0000000000;
	notes[371] = 10'b0010000100;
	notes[372] = 10'b0001000010;
	notes[373] = 10'b0000000000;
	notes[374] = 10'b0001000010;
	notes[375] = 10'b0000000000;
	notes[376] = 10'b1000001010; // 50
	notes[377] = 10'b0000000000;
	notes[378] = 10'b0000000000;
	notes[379] = 10'b1000001010;
	notes[380] = 10'b1000001010;
	notes[381] = 10'b0000000000;
	notes[382] = 10'b0000000000;
	notes[383] = 10'b0000000000;
	notes[384] = 10'b0010001100; // 51
	notes[385] = 10'b0010001100;
	notes[386] = 10'b0000000000;
	notes[387] = 10'b0010000100;
	notes[388] = 10'b0001000010;
	notes[389] = 10'b0000000000;
	notes[390] = 10'b0001000010;
	notes[391] = 10'b0000000000;
	notes[392] = 10'b0100010100; // 52
	notes[393] = 10'b0100010100;
	notes[394] = 10'b0000000000;
	notes[395] = 10'b0100010100;
	notes[396] = 10'b0100010100;
	notes[397] = 10'b0100010100;
	notes[398] = 10'b0000000000;
	notes[399] = 10'b0100010100;
	notes[400] = 10'b0010001100; // 53
	notes[401] = 10'b0010001100;
	notes[402] = 10'b0000000000;
	notes[403] = 10'b0010000100;
	notes[404] = 10'b0001000010;
	notes[405] = 10'b0000000000;
	notes[406] = 10'b0001000010;
	notes[407] = 10'b0000000000;
	notes[408] = 10'b1000011000; // 54
	notes[409] = 10'b1000011000;
	notes[410] = 10'b0000000000;
	notes[411] = 10'b1000011000;
	notes[412] = 10'b1000011000;
	notes[413] = 10'b1000011000;
	notes[414] = 10'b0000000000;
	notes[415] = 10'b0000011000;
	notes[416] = 10'b0010001100; // 55
	notes[417] = 10'b0010001100;
	notes[418] = 10'b0000000000;
	notes[419] = 10'b0010000100;
	notes[420] = 10'b0001000010;
	notes[421] = 10'b0000000000;
	notes[422] = 10'b0001000010;
	notes[423] = 10'b0000000000;
	notes[424] = 10'b0100010100; // 56
	notes[425] = 10'b0100010100;
	notes[426] = 10'b0000000000;
	notes[427] = 10'b0100010100;
	notes[428] = 10'b0100010100;
	notes[429] = 10'b0100010100;
	notes[430] = 10'b0000000000;
	notes[431] = 10'b0100010100;
	notes[432] = 10'b0010001100; // 57
	notes[433] = 10'b0010001100;
	notes[434] = 10'b0000000000;
	notes[435] = 10'b0010000100;
	notes[436] = 10'b0001000010;
	notes[437] = 10'b0000000000;
	notes[438] = 10'b0001000010;
	notes[439] = 10'b0000000000;
	notes[440] = 10'b0010001010; // 58
	notes[441] = 10'b0010001010;
	notes[442] = 10'b0010001010;
	notes[443] = 10'b0010000000;
	notes[444] = 10'b0100001100;
	notes[445] = 10'b0100001100;
	notes[446] = 10'b0100001100;
	notes[447] = 10'b0100000000;
	notes[448] = 10'b0010001000; // 59
	notes[449] = 10'b0010000000;
	notes[450] = 10'b0000001000;
	notes[451] = 10'b0010001000;
	notes[452] = 10'b0001001000;
	notes[453] = 10'b0000000100;
	notes[454] = 10'b0001001000;
	notes[455] = 10'b0000000100;
	notes[456] = 10'b0100001000; // 60
	notes[457] = 10'b0100000000;
	notes[458] = 10'b0000001000;
	notes[459] = 10'b0100001000;
	notes[460] = 10'b0100001000;
	notes[461] = 10'b0100000100;
	notes[462] = 10'b0000001000;
	notes[463] = 10'b0100000100;
	notes[464] = 10'b0010001000; // 61
	notes[465] = 10'b0010000000;
	notes[466] = 10'b0000001000;
	notes[467] = 10'b0010001000;
	notes[468] = 10'b0001001000;
	notes[469] = 10'b0000000100;
	notes[470] = 10'b0001001000;
	notes[471] = 10'b0000000100;
	notes[472] = 10'b1000001000; // 62
	notes[473] = 10'b1000000000;
	notes[474] = 10'b0000001000;
	notes[475] = 10'b1000001000;
	notes[476] = 10'b1000001000;
	notes[477] = 10'b1000010000;
	notes[478] = 10'b0000010000;
	notes[479] = 10'b0000010000;
	notes[480] = 10'b0010001000; // 63
	notes[481] = 10'b0010000000;
	notes[482] = 10'b0000001000;
	notes[483] = 10'b0010001000;
	notes[484] = 10'b0001001000;
	notes[485] = 10'b0000000100;
	notes[486] = 10'b0001001000;
	notes[487] = 10'b0000000100;
	notes[488] = 10'b0100001000; // 64
	notes[489] = 10'b0100000000;
	notes[490] = 10'b0000001000;
	notes[491] = 10'b0100001000;
	notes[492] = 10'b0100001000;
	notes[493] = 10'b0100000100;
	notes[494] = 10'b0000001000;
	notes[495] = 10'b0100000100;
	notes[496] = 10'b0010001000; // 65
	notes[497] = 10'b0010000000;
	notes[498] = 10'b0000001000;
	notes[499] = 10'b0010001000;
	notes[500] = 10'b0001001000;
	notes[501] = 10'b0000000100;
	notes[502] = 10'b0001001000;
	notes[503] = 10'b0000000100;
	notes[504] = 10'b0010000010; // 66
	notes[505] = 10'b0010000000;
	notes[506] = 10'b0010000010;
	notes[507] = 10'b0010000010;
	notes[508] = 10'b0100000010;
	notes[509] = 10'b0100000001;
	notes[510] = 10'b0100000001;
	notes[511] = 10'b0100000000;
	notes[512] = 10'b0001001010; // 67
	notes[513] = 10'b0001001010;
	notes[514] = 10'b0001001010;
	notes[515] = 10'b0001001010;
	notes[516] = 10'b0001001010;
	notes[517] = 10'b0001001010;
	notes[518] = 10'b0001001010;
	notes[519] = 10'b0001000000;
	notes[520] = 10'b0100010100; // 68
	notes[521] = 10'b0100010100;
	notes[522] = 10'b0100010100;
	notes[523] = 10'b0100010100;
	notes[524] = 10'b0100010100;
	notes[525] = 10'b0000000000;
	notes[526] = 10'b0000000000;
	notes[527] = 10'b0000000000;
	notes[528] = 10'b1000001010; // 69
	notes[529] = 10'b0000000000;
	notes[530] = 10'b1000001010;
	notes[531] = 10'b0000000000;
	notes[532] = 10'b0001001010;
	notes[533] = 10'b0000100000;
	notes[534] = 10'b0001001010;
	notes[535] = 10'b0000000000;
	notes[536] = 10'b0010001100; // 70
	notes[537] = 10'b0000000000;
	notes[538] = 10'b0010001100;
	notes[539] = 10'b0000000000;
	notes[540] = 10'b0010001100;
	notes[541] = 10'b0000100000;
	notes[542] = 10'b0010001100;
	notes[543] = 10'b0000000000;
	notes[544] = 10'b1000010010; // 71
	notes[545] = 10'b0000000000;
	notes[546] = 10'b1000010010;
	notes[547] = 10'b0000000000;
	notes[548] = 10'b1000010010;
	notes[549] = 10'b0010000000;
	notes[550] = 10'b1000010010;
	notes[551] = 10'b0000000000;
	notes[552] = 10'b0100000101; // 72
	notes[553] = 10'b0100000000;
	notes[554] = 10'b0100000101;
	notes[555] = 10'b0100000000;
	notes[556] = 10'b0010000110;
	notes[557] = 10'b0010000000;
	notes[558] = 10'b0010000110;
	notes[559] = 10'b0010000000;
	notes[560] = 10'b0001001010; // 73
	notes[561] = 10'b0000000000;
	notes[562] = 10'b0001001010;
	notes[563] = 10'b0000000000;
	notes[564] = 10'b0001001010;
	notes[565] = 10'b0000100000;
	notes[566] = 10'b0001001010;
	notes[567] = 10'b0000000000;
	notes[568] = 10'b0010001100; // 74
	notes[569] = 10'b0000000000;
	notes[570] = 10'b0010001100;
	notes[571] = 10'b0000000000;
	notes[572] = 10'b0010001100;
	notes[573] = 10'b0001000000;
	notes[574] = 10'b0010001100;
	notes[575] = 10'b0000000000;
	notes[576] = 10'b1000010010; // 75
	notes[577] = 10'b0000000000;
	notes[578] = 10'b1000010010;
	notes[579] = 10'b0000000000;
	notes[580] = 10'b1000010010;
	notes[581] = 10'b0010000000;
	notes[582] = 10'b1000010010;
	notes[583] = 10'b0000000000;
	notes[584] = 10'b0100000101; // 76
	notes[585] = 10'b0100000000;
	notes[586] = 10'b0100000101;
	notes[587] = 10'b0100000000;
	notes[588] = 10'b0010000110;
	notes[589] = 10'b0010000000;
	notes[590] = 10'b0010000110;
	notes[591] = 10'b0010000000;
	notes[592] = 10'b0001001010; // 77
	notes[593] = 10'b0000000000;
	notes[594] = 10'b0001001010;
	notes[595] = 10'b0000000000;
	notes[596] = 10'b0001001010;
	notes[597] = 10'b0000000000;
	notes[598] = 10'b0001001010;
	notes[599] = 10'b0000000000;
	notes[600] = 10'b0001001010; // 78
	notes[601] = 10'b0000000000;
	notes[602] = 10'b0001001010;
	notes[603] = 10'b0000000000;
	notes[604] = 10'b0001001010;
	notes[605] = 10'b0010000101;
	notes[606] = 10'b0010000101;
	notes[607] = 10'b0010000000;
	notes[608] = 10'b1000000110; // 79
	notes[609] = 10'b0000000000;
	notes[610] = 10'b1000000110;
	notes[611] = 10'b0000000000;
	notes[612] = 10'b1000000110;
	notes[613] = 10'b0000000000;
	notes[614] = 10'b1000000110;
	notes[615] = 10'b0000000000;
	notes[616] = 10'b1000000110; // 80
	notes[617] = 10'b0000000000;
	notes[618] = 10'b1000000110;
	notes[619] = 10'b0000000000;
	notes[620] = 10'b1000000110;
	notes[621] = 10'b0100000101;
	notes[622] = 10'b0100000101;
	notes[623] = 10'b0010000000;
	notes[624] = 10'b0001001010; // 81
	notes[625] = 10'b0000000000;
	notes[626] = 10'b0001001010;
	notes[627] = 10'b0000000000;
	notes[628] = 10'b0001001010;
	notes[629] = 10'b0000000000;
	notes[630] = 10'b0001001010;
	notes[631] = 10'b0000000000;
	notes[632] = 10'b0001001010; // 82
	notes[633] = 10'b0000000000;
	notes[634] = 10'b0001001010;
	notes[635] = 10'b0000000000;
	notes[636] = 10'b0001001010;
	notes[637] = 10'b0010000101;
	notes[638] = 10'b0010000101;
	notes[639] = 10'b0010000000;
	notes[640] = 10'b1000000110; // 83
	notes[641] = 10'b0000000000;
	notes[642] = 10'b1000000110;
	notes[643] = 10'b0000000000;
	notes[644] = 10'b1000000110;
	notes[645] = 10'b0000000000;
	notes[646] = 10'b1000000110;
	notes[647] = 10'b0000000000;
	notes[648] = 10'b0010000001; // 84
	notes[649] = 10'b0010000001;
	notes[650] = 10'b0010000001;
	notes[651] = 10'b0010000001;
	notes[652] = 10'b0100000010;
	notes[653] = 10'b0000000000;
	notes[654] = 10'b0000000000;
	notes[655] = 10'b0000000000;
	notes[656] = 10'b0000000011; // 85
	notes[657] = 10'b0000000000;
	notes[658] = 10'b0000000100;
	notes[659] = 10'b0000000001;
	notes[660] = 10'b0000000000;
	notes[661] = 10'b0000000000;
	notes[662] = 10'b0000000100;
	notes[663] = 10'b0000000000;
	notes[664] = 10'b0000000101; // 86
	notes[665] = 10'b0000000000;
	notes[666] = 10'b0000000100;
	notes[667] = 10'b0000000001;
	notes[668] = 10'b0000000000;
	notes[669] = 10'b0000000000;
	notes[670] = 10'b0000001000;
	notes[671] = 10'b0000000000;
	notes[672] = 10'b0000001010; // 87
	notes[673] = 10'b0000000000;
	notes[674] = 10'b0000001000;
	notes[675] = 10'b0000000001;
	notes[676] = 10'b0000000000;
	notes[677] = 10'b0000000000;
	notes[678] = 10'b0000001000;
	notes[679] = 10'b0000000000;
	notes[680] = 10'b0000001010; // 88
	notes[681] = 10'b0000000000;
	notes[682] = 10'b0000000000;
	notes[683] = 10'b0000000000;
	notes[684] = 10'b0000010010;
	notes[685] = 10'b0000000000;
	notes[686] = 10'b0000000000;
	notes[687] = 10'b0000000000;
	notes[688] = 10'b0010000011; // 89
	notes[689] = 10'b0000000000;
	notes[690] = 10'b0000000100;
	notes[691] = 10'b0000000001;
	notes[692] = 10'b0000000000;
	notes[693] = 10'b0000000000;
	notes[694] = 10'b0010000100;
	notes[695] = 10'b0000000000;
	notes[696] = 10'b0000100101; // 90
	notes[697] = 10'b0000000000;
	notes[698] = 10'b0000000100;
	notes[699] = 10'b0000000001;
	notes[700] = 10'b0000000000;
	notes[701] = 10'b0000000000;
	notes[702] = 10'b0000001000;
	notes[703] = 10'b0000000000;
	notes[704] = 10'b0100001010; // 91
	notes[705] = 10'b0000000000;
	notes[706] = 10'b0000001000;
	notes[707] = 10'b0000000001;
	notes[708] = 10'b0000000000;
	notes[709] = 10'b0000000000;
	notes[710] = 10'b0000001000;
	notes[711] = 10'b0000000000;
	notes[712] = 10'b0010001010; // 92
	notes[713] = 10'b0000000000;
	notes[714] = 10'b0000000000;
	notes[715] = 10'b0000000000;
	notes[716] = 10'b0001010010;
	notes[717] = 10'b0000000000;
	notes[718] = 10'b0000000000;
	notes[719] = 10'b0000000000;
	notes[720] = 10'b0010000011; // 93
	notes[721] = 10'b0000000000;
	notes[722] = 10'b0000000100;
	notes[723] = 10'b0000000001;
	notes[724] = 10'b0000000000;
	notes[725] = 10'b0000000000;
	notes[726] = 10'b0000000100;
	notes[727] = 10'b0000000000;
	notes[728] = 10'b0100000101; // 94
	notes[729] = 10'b0000000000;
	notes[730] = 10'b0000000100;
	notes[731] = 10'b0000000001;
	notes[732] = 10'b0000000000;
	notes[733] = 10'b0000000000;
	notes[734] = 10'b0000001000;
	notes[735] = 10'b0000000000;
	notes[736] = 10'b1000001010; // 95
	notes[737] = 10'b0000000000;
	notes[738] = 10'b0000001000;
	notes[739] = 10'b0000000001;
	notes[740] = 10'b0000000000;
	notes[741] = 10'b0000000000;
	notes[742] = 10'b0000001000;
	notes[743] = 10'b0000000000;
	notes[744] = 10'b0010001010; // 96
	notes[745] = 10'b0000000000;
	notes[746] = 10'b0000000000;
	notes[747] = 10'b0000000000;
	notes[748] = 10'b0001010010;
	notes[749] = 10'b0000000000;
	notes[750] = 10'b0000000000;
	notes[751] = 10'b0000000000;
	notes[752] = 10'b0010000011; // 97
	notes[753] = 10'b0000000000;
	notes[754] = 10'b0000000100;
	notes[755] = 10'b0000000001;
	notes[756] = 10'b0000000000;
	notes[757] = 10'b0000000000;
	notes[758] = 10'b0010000100;
	notes[759] = 10'b0000000000;
	notes[760] = 10'b0000100101; // 98
	notes[761] = 10'b0000000000;
	notes[762] = 10'b0000000100;
	notes[763] = 10'b0000000001;
	notes[764] = 10'b0000000000;
	notes[765] = 10'b0000000000;
	notes[766] = 10'b0000001000;
	notes[767] = 10'b0000000000;
	notes[768] = 10'b0100001010; // 99
	notes[769] = 10'b0000000000;
	notes[770] = 10'b0000001000;
	notes[771] = 10'b0000000001;
	notes[772] = 10'b0000000000;
	notes[773] = 10'b0000000000;
	notes[774] = 10'b0000001000;
	notes[775] = 10'b0000000000;
	notes[776] = 10'b0010001010; // 100
	notes[777] = 10'b0010000000;
	notes[778] = 10'b0010000000;
	notes[779] = 10'b0010000000;
	notes[780] = 10'b0010010010;
	notes[781] = 10'b0000000000;
	notes[782] = 10'b0000000000;
	notes[783] = 10'b0000000000;
	notes[784] = 10'b0001010000; // 101
	notes[785] = 10'b0000001000;
	notes[786] = 10'b0001001000;
	notes[787] = 10'b0000001000;
	notes[788] = 10'b0001001000;
	notes[789] = 10'b0000101000;
	notes[790] = 10'b0001001000;
	notes[791] = 10'b0000000000;
	notes[792] = 10'b0010010000; // 102
	notes[793] = 10'b0000001000;
	notes[794] = 10'b0010001000;
	notes[795] = 10'b0000001000;
	notes[796] = 10'b0010001000;
	notes[797] = 10'b0000101000;
	notes[798] = 10'b0010001000;
	notes[799] = 10'b0000000000;
	notes[800] = 10'b1000010000; // 103
	notes[801] = 10'b0000001000;
	notes[802] = 10'b1000001000;
	notes[803] = 10'b0000001000;
	notes[804] = 10'b1000001000;
	notes[805] = 10'b0010001000;
	notes[806] = 10'b1000001000;
	notes[807] = 10'b0000000000;
	notes[808] = 10'b0100000001; // 104
	notes[809] = 10'b0100000001;
	notes[810] = 10'b0100000001;
	notes[811] = 10'b0100000000;
	notes[812] = 10'b0010000100;
	notes[813] = 10'b0010000100;
	notes[814] = 10'b0010000100;
	notes[815] = 10'b0010000000;
	notes[816] = 10'b0001010000; // 105
	notes[817] = 10'b0000001000;
	notes[818] = 10'b0001001000;
	notes[819] = 10'b0000001000;
	notes[820] = 10'b0001001000;
	notes[821] = 10'b0000101000;
	notes[822] = 10'b0001001000;
	notes[823] = 10'b0000000000;
	notes[824] = 10'b0100010000; // 106
	notes[825] = 10'b0000001000;
	notes[826] = 10'b0100001000;
	notes[827] = 10'b0000001000;
	notes[828] = 10'b0100001000;
	notes[829] = 10'b0010001000;
	notes[830] = 10'b0100001000;
	notes[831] = 10'b0000000000;
	notes[832] = 10'b1000010000; // 107
	notes[833] = 10'b0000001000;
	notes[834] = 10'b1000001000;
	notes[835] = 10'b0000001000;
	notes[836] = 10'b1000001000;
	notes[837] = 10'b0100001000;
	notes[838] = 10'b1000001000;
	notes[839] = 10'b0000000000;
	notes[840] = 10'b0100000001; // 108
	notes[841] = 10'b0100000001;
	notes[842] = 10'b0100000001;
	notes[843] = 10'b0100000000;
	notes[844] = 10'b0010000100;
	notes[845] = 10'b0010000100;
	notes[846] = 10'b0010000100;
	notes[847] = 10'b0010000000;
	notes[848] = 10'b0001000010; // 109
	notes[849] = 10'b0001000010;
	notes[850] = 10'b0001000010;
	notes[851] = 10'b0001000010;
	notes[852] = 10'b0001000010;
	notes[853] = 10'b0001000010;
	notes[854] = 10'b0001000010;
	notes[855] = 10'b0001000000;
	notes[856] = 10'b0001000100; // 110
	notes[857] = 10'b0001000100;
	notes[858] = 10'b0001000100;
	notes[859] = 10'b0001000100;
	notes[860] = 10'b0001000100;
	notes[861] = 10'b0010000100;
	notes[862] = 10'b0010000100;
	notes[863] = 10'b0010000000;
	notes[864] = 10'b1000001000; // 111
	notes[865] = 10'b1000001000;
	notes[866] = 10'b1000001000;
	notes[867] = 10'b1000001000;
	notes[868] = 10'b1000001000;
	notes[869] = 10'b1000001000;
	notes[870] = 10'b1000001000;
	notes[871] = 10'b1000000000;
	notes[872] = 10'b1000010000; // 112
	notes[873] = 10'b1000010000;
	notes[874] = 10'b1000010000;
	notes[875] = 10'b1000010000;
	notes[876] = 10'b1000010000;
	notes[877] = 10'b0100010000;
	notes[878] = 10'b0100010000;
	notes[879] = 10'b0100000000;
	notes[880] = 10'b0001000010; // 113
	notes[881] = 10'b0001000010;
	notes[882] = 10'b0001000010;
	notes[883] = 10'b0001000010;
	notes[884] = 10'b0001000010;
	notes[885] = 10'b0001000010;
	notes[886] = 10'b0001000010;
	notes[887] = 10'b0001000000;
	notes[888] = 10'b0001000001; // 114
	notes[889] = 10'b0001000001;
	notes[890] = 10'b0001000001;
	notes[891] = 10'b0001000001;
	notes[892] = 10'b0001000001;
	notes[893] = 10'b0010000001;
	notes[894] = 10'b0010000001;
	notes[895] = 10'b0010000000;
	notes[896] = 10'b1000000100; // 115
	notes[897] = 10'b1000000100;
	notes[898] = 10'b1000000100;
	notes[899] = 10'b1000000000;
	notes[900] = 10'b1000000010;
	notes[901] = 10'b1000000010;
	notes[902] = 10'b1000000001;
	notes[903] = 10'b1000000000;
	notes[904] = 10'b0010000010; // 116
	notes[905] = 10'b0010000010;
	notes[906] = 10'b0010000010;
	notes[907] = 10'b0010000000;
	notes[908] = 10'b0100000010;
	notes[909] = 10'b0000000000;
	notes[910] = 10'b0000000000;
	notes[911] = 10'b0000000000;
	notes[912] = 10'b0000000000; // 117
	notes[913] = 10'b0000000000;
	notes[914] = 10'b0000000000;
	notes[915] = 10'b0000000000;
	notes[916] = 10'b0000000000;
	notes[917] = 10'b0000000000;
	notes[918] = 10'b0000000000;
	notes[919] = 10'b0000000000;
	notes[920] = 10'b0000000000; // 118
	notes[921] = 10'b0000000000;
	notes[922] = 10'b0000000000;
	notes[923] = 10'b0000000000;
	notes[924] = 10'b0000000000;
	notes[925] = 10'b0000000000;
	notes[926] = 10'b0000000000;
	notes[927] = 10'b0000000000;
	notes[928] = 10'b0000000000; // 119
	notes[929] = 10'b0000000000;
	notes[930] = 10'b0000000000;
	notes[931] = 10'b0000000000;
	notes[932] = 10'b0000000000;
	notes[933] = 10'b0000000000;
	notes[934] = 10'b0000000000;
	notes[935] = 10'b0000000000;
	notes[936] = 10'b0000000000; // 120
	notes[937] = 10'b0000000000;
	notes[938] = 10'b0000000000;
	notes[939] = 10'b0000000000;
	notes[940] = 10'b0000000000;
	notes[941] = 10'b0000000000;
	notes[942] = 10'b0000000000;
	notes[943] = 10'b0000000000;
	notes[944] = 10'b1000001010; // 121
	notes[945] = 10'b0000000000;
	notes[946] = 10'b1000001010;
	notes[947] = 10'b0000000000;
	notes[948] = 10'b1000001010;
	notes[949] = 10'b0100000000;
	notes[950] = 10'b1000001010;
	notes[951] = 10'b1000000000;
	notes[952] = 10'b0010001100; // 122
	notes[953] = 10'b0000000000;
	notes[954] = 10'b0010001100;
	notes[955] = 10'b0000000000;
	notes[956] = 10'b0010001100;
	notes[957] = 10'b0001000000;
	notes[958] = 10'b0010001100;
	notes[959] = 10'b0000000000;
	notes[960] = 10'b1000010010; // 123
	notes[961] = 10'b0000000000;
	notes[962] = 10'b1000010010;
	notes[963] = 10'b0000000000;
	notes[964] = 10'b1000010010;
	notes[965] = 10'b0100000000;
	notes[966] = 10'b1000010010;
	notes[967] = 10'b0000000000;
	notes[968] = 10'b0100000101; // 124
	notes[969] = 10'b0100000000;
	notes[970] = 10'b0100000101;
	notes[971] = 10'b0100000000;
	notes[972] = 10'b0010000110;
	notes[973] = 10'b0010000000;
	notes[974] = 10'b0010000110;
	notes[975] = 10'b0010000000;
	notes[976] = 10'b0001001010; // 125
	notes[977] = 10'b0000000000;
	notes[978] = 10'b0001001010;
	notes[979] = 10'b0000000000;
	notes[980] = 10'b0001001010;
	notes[981] = 10'b0000100000;
	notes[982] = 10'b0001001010;
	notes[983] = 10'b0000000000;
	notes[984] = 10'b0100001100; // 126
	notes[985] = 10'b0000000000;
	notes[986] = 10'b0100001100;
	notes[987] = 10'b0000000000;
	notes[988] = 10'b0100001100;
	notes[989] = 10'b0010000000;
	notes[990] = 10'b0100001100;
	notes[991] = 10'b0000000000;
	notes[992] = 10'b1000010010; // 127
	notes[993] = 10'b0000000000;
	notes[994] = 10'b1000010010;
	notes[995] = 10'b0000000000;
	notes[996] = 10'b1000010010;
	notes[997] = 10'b0010000000;
	notes[998] = 10'b1000010010;
	notes[999] = 10'b0000000000;
	notes[1000] = 10'b0100000101; // 128
	notes[1001] = 10'b0100000000;
	notes[1002] = 10'b0100000101;
	notes[1003] = 10'b0100000000;
	notes[1004] = 10'b0010000110;
	notes[1005] = 10'b0010000000;
	notes[1006] = 10'b0010000110;
	notes[1007] = 10'b0010000000;
	notes[1008] = 10'b0001001010; // 129
	notes[1009] = 10'b0000000000;
	notes[1010] = 10'b0001001010;
	notes[1011] = 10'b0000000000;
	notes[1012] = 10'b0001001010;
	notes[1013] = 10'b0000000000;
	notes[1014] = 10'b0001001010;
	notes[1015] = 10'b0000000000;
	notes[1016] = 10'b0001001010; // 130
	notes[1017] = 10'b0000000000;
	notes[1018] = 10'b0001001010;
	notes[1019] = 10'b0000000000;
	notes[1020] = 10'b0001001010;
	notes[1021] = 10'b0010000101;
	notes[1022] = 10'b0010000101;
	notes[1023] = 10'b0010000000;
	notes[1024] = 10'b1000000110; // 131
	notes[1025] = 10'b0000000000;
	notes[1026] = 10'b1000000110;
	notes[1027] = 10'b0000000000;
	notes[1028] = 10'b1000000110;
	notes[1029] = 10'b0000000000;
	notes[1030] = 10'b1000000110;
	notes[1031] = 10'b0000000000;
	notes[1032] = 10'b1000000110; // 132
	notes[1033] = 10'b0000000000;
	notes[1034] = 10'b1000000110;
	notes[1035] = 10'b0000000000;
	notes[1036] = 10'b1000000110;
	notes[1037] = 10'b0100000101;
	notes[1038] = 10'b0100000101;
	notes[1039] = 10'b0010000000;
	notes[1040] = 10'b0001001010; // 133
	notes[1041] = 10'b0000000000;
	notes[1042] = 10'b0001001010;
	notes[1043] = 10'b0000000000;
	notes[1044] = 10'b0001001010;
	notes[1045] = 10'b0000000000;
	notes[1046] = 10'b0001001010;
	notes[1047] = 10'b0000000000;
	notes[1048] = 10'b0001001010; // 134
	notes[1049] = 10'b0000000000;
	notes[1050] = 10'b0001001010;
	notes[1051] = 10'b0000000000;
	notes[1052] = 10'b0001001010;
	notes[1053] = 10'b0010000101;
	notes[1054] = 10'b0010000101;
	notes[1055] = 10'b0010000000;
	notes[1056] = 10'b1000000110; // 135
	notes[1057] = 10'b0000000000;
	notes[1058] = 10'b1000000110;
	notes[1059] = 10'b0000000000;
	notes[1060] = 10'b1000000110;
	notes[1061] = 10'b0000000000;
	notes[1062] = 10'b1000000110;
	notes[1063] = 10'b0000000000;
	notes[1064] = 10'b0010000001; // 136
	notes[1065] = 10'b0010000001;
	notes[1066] = 10'b0010000001;
	notes[1067] = 10'b0010000001;
	notes[1068] = 10'b0100000010;
	notes[1069] = 10'b0000000000;
	notes[1070] = 10'b0000000000;
	notes[1071] = 10'b0000000000;
	notes[1072] = 10'b0010000100; // 137
	notes[1073] = 10'b0010000100;
	notes[1074] = 10'b0000000000;
	notes[1075] = 10'b0010000100;
	notes[1076] = 10'b0001000010;
	notes[1077] = 10'b0000000000;
	notes[1078] = 10'b0001000010;
	notes[1079] = 10'b0000000000;
	notes[1080] = 10'b0100001000; // 138
	notes[1081] = 10'b0100001000;
	notes[1082] = 10'b0000000000;
	notes[1083] = 10'b0100001000;
	notes[1084] = 10'b0100001000;
	notes[1085] = 10'b0100001000;
	notes[1086] = 10'b0000000000;
	notes[1087] = 10'b0100001000;
	notes[1088] = 10'b0010000100; // 139
	notes[1089] = 10'b0010000100;
	notes[1090] = 10'b0000000000;
	notes[1091] = 10'b0010000100;
	notes[1092] = 10'b0001000010;
	notes[1093] = 10'b0000000000;
	notes[1094] = 10'b0001000010;
	notes[1095] = 10'b0000000000;
	notes[1096] = 10'b1000010000; // 140
	notes[1097] = 10'b1000010000;
	notes[1098] = 10'b0000000000;
	notes[1099] = 10'b1000010000;
	notes[1100] = 10'b1000010000;
	notes[1101] = 10'b1000010000;
	notes[1102] = 10'b0000000000;
	notes[1103] = 10'b0000000000;
	notes[1104] = 10'b0010000100; // 141
	notes[1105] = 10'b0010000100;
	notes[1106] = 10'b0000000000;
	notes[1107] = 10'b0010000100;
	notes[1108] = 10'b0001000010;
	notes[1109] = 10'b0000000000;
	notes[1110] = 10'b0001000010;
	notes[1111] = 10'b0000000000;
	notes[1112] = 10'b0100001000; // 142
	notes[1113] = 10'b0100001000;
	notes[1114] = 10'b0000000000;
	notes[1115] = 10'b0100001000;
	notes[1116] = 10'b0100001000;
	notes[1117] = 10'b0100001000;
	notes[1118] = 10'b0000000000;
	notes[1119] = 10'b0100001000;
	notes[1120] = 10'b0010000100; // 143
	notes[1121] = 10'b0010000100;
	notes[1122] = 10'b0000000000;
	notes[1123] = 10'b0010000100;
	notes[1124] = 10'b0001000010;
	notes[1125] = 10'b0000000000;
	notes[1126] = 10'b0000000000;
	notes[1127] = 10'b0000000000;
	notes[1128] = 10'b1000010000; // 144
	notes[1129] = 10'b0000000000;
	notes[1130] = 10'b0000000000;
	notes[1131] = 10'b1000010000;
	notes[1132] = 10'b1000010000;
	notes[1133] = 10'b0000000000;
	notes[1134] = 10'b0000000000;
	notes[1135] = 10'b0000000000;
	notes[1136] = 10'b0000000000; // fin.
	notes[1137] = 10'b0000000000;
	notes[1138] = 10'b0000000000;
	notes[1139] = 10'b0000000000;
	notes[1140] = 10'b0000000000;
	notes[1141] = 10'b0000000000;
	notes[1142] = 10'b0000000000;
	notes[1143] = 10'b0000000000;
	notes[1144] = 10'b0000000000;
	notes[1145] = 10'b0000000000;
	notes[1146] = 10'b0000000000;
	notes[1147] = 10'b0000000000;
	notes[1148] = 10'b0000000000;
	notes[1149] = 10'b0000000000;
	notes[1150] = 10'b0000000000;
	notes[1151] = 10'b0000000000;
	notes[1152] = 10'b0000000000;
	notes[1153] = 10'b0000000000;
	notes[1154] = 10'b0000000000;
	notes[1155] = 10'b0000000000;
	notes[1156] = 10'b0000000000;
	notes[1157] = 10'b0000000000;
	notes[1158] = 10'b0000000000;
	notes[1159] = 10'b0000000000;
	notes[1160] = 10'b0000000000;
	notes[1161] = 10'b0000000000;
	notes[1162] = 10'b0000000000;
	notes[1163] = 10'b0000000000;
	notes[1164] = 10'b0000000000;
	notes[1165] = 10'b0000000000;
	notes[1166] = 10'b0000000000;
	notes[1167] = 10'b0000000000;
	notes[1168] = 10'b0000000000;
	notes[1169] = 10'b0000000000;
	notes[1170] = 10'b0000000000;
	notes[1171] = 10'b0000000000;
	notes[1172] = 10'b0000000000;
	notes[1173] = 10'b0000000000;
	notes[1174] = 10'b0000000000;
	notes[1175] = 10'b0000000000;
	notes[1176] = 10'b0000000000;
	notes[1177] = 10'b0000000000;
	notes[1178] = 10'b0000000000;
	notes[1179] = 10'b0000000000;
	notes[1180] = 10'b0000000000;
	notes[1181] = 10'b0000000000;
	notes[1182] = 10'b0000000000;
	notes[1183] = 10'b0000000000;
	notes[1184] = 10'b0000000000;
	notes[1185] = 10'b0000000000;
	notes[1186] = 10'b0000000000;
	notes[1187] = 10'b0000000000;
	notes[1188] = 10'b0000000000;
	notes[1189] = 10'b0000000000;
	notes[1190] = 10'b0000000000;
	notes[1191] = 10'b0000000000;
	notes[1192] = 10'b0000000000;
	notes[1193] = 10'b0000000000;
	notes[1194] = 10'b0000000000;
	notes[1195] = 10'b0000000000;
	notes[1196] = 10'b0000000000;
	notes[1197] = 10'b0000000000;
	notes[1198] = 10'b0000000000;
	notes[1199] = 10'b0000000000;

end

always_ff @(posedge clk) begin
	data <= notes[addr];
end

endmodule
